module leds_on(output wire [7:0] LPORT);

//-- Turn on all the leds
assign LPORT = 8'hFF;

endmodule
